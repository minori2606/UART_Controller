library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity mFlashMem is
	Port (
		adr : in  STD_LOGIC_VECTOR (15 downto 0);
		dat : out  STD_LOGIC_VECTOR (15 downto 0));
end mFlashMem;

architecture Behavioral of mFlashMem is

begin
	process (adr) begin
		case (adr) is
			when x"0000" => dat <= x"120A";
			when x"0001" => dat <= x"118A";
			when x"0002" => dat <= x"2803";
			when x"0003" => dat <= x"1003";
			when x"0004" => dat <= x"3000";
			when x"0005" => dat <= x"1803";
			when x"0006" => dat <= x"3001";
			when x"0007" => dat <= x"00A4";
			when x"0008" => dat <= x"1003";
			when x"0009" => dat <= x"3000";
			when x"000A" => dat <= x"1803";
			when x"000B" => dat <= x"3001";
			when x"000C" => dat <= x"00A6";
			when x"000D" => dat <= x"3000";
			when x"000E" => dat <= x"1283";
			when x"000F" => dat <= x"1703";
			when x"0010" => dat <= x"0093";
			when x"0011" => dat <= x"3000";
			when x"0012" => dat <= x"0094";
			when x"0013" => dat <= x"2814";
			when x"0014" => dat <= x"1003";
			when x"0015" => dat <= x"0813";
			when x"0016" => dat <= x"3E15";
			when x"0017" => dat <= x"1783";
			when x"0018" => dat <= x"0084";
			when x"0019" => dat <= x"3000";
			when x"001A" => dat <= x"1803";
			when x"001B" => dat <= x"3001";
			when x"001C" => dat <= x"0080";
			when x"001D" => dat <= x"3001";
			when x"001E" => dat <= x"0793";
			when x"001F" => dat <= x"1803";
			when x"0020" => dat <= x"0A94";
			when x"0021" => dat <= x"3000";
			when x"0022" => dat <= x"0794";
			when x"0023" => dat <= x"0814";
			when x"0024" => dat <= x"3A80";
			when x"0025" => dat <= x"00D5";
			when x"0026" => dat <= x"3080";
			when x"0027" => dat <= x"0255";
			when x"0028" => dat <= x"1D03";
			when x"0029" => dat <= x"282C";
			when x"002A" => dat <= x"3040";
			when x"002B" => dat <= x"0213";
			when x"002C" => dat <= x"1C03";
			when x"002D" => dat <= x"282F";
			when x"002E" => dat <= x"2830";
			when x"002F" => dat <= x"2814";
			when x"0030" => dat <= x"1283";
			when x"0031" => dat <= x"1303";
			when x"0032" => dat <= x"0823";
			when x"0033" => dat <= x"3920";
			when x"0034" => dat <= x"1283";
			when x"0035" => dat <= x"1703";
			when x"0036" => dat <= x"0090";
			when x"0037" => dat <= x"0810";
			when x"0038" => dat <= x"3A20";
			when x"0039" => dat <= x"1D03";
			when x"003A" => dat <= x"283C";
			when x"003B" => dat <= x"283D";
			when x"003C" => dat <= x"2899";
			when x"003D" => dat <= x"3015";
			when x"003E" => dat <= x"120A";
			when x"003F" => dat <= x"118A";
			when x"0040" => dat <= x"2720";
			when x"0041" => dat <= x"120A";
			when x"0042" => dat <= x"118A";
			when x"0043" => dat <= x"1283";
			when x"0044" => dat <= x"1703";
			when x"0045" => dat <= x"0857";
			when x"0046" => dat <= x"0194";
			when x"0047" => dat <= x"0794";
			when x"0048" => dat <= x"0856";
			when x"0049" => dat <= x"0193";
			when x"004A" => dat <= x"0793";
			when x"004B" => dat <= x"3000";
			when x"004C" => dat <= x"0091";
			when x"004D" => dat <= x"3000";
			when x"004E" => dat <= x"0092";
			when x"004F" => dat <= x"2872";
			when x"0050" => dat <= x"3001";
			when x"0051" => dat <= x"00D5";
			when x"0052" => dat <= x"1283";
			when x"0053" => dat <= x"1303";
			when x"0054" => dat <= x"1283";
			when x"0055" => dat <= x"1703";
			when x"0056" => dat <= x"0855";
			when x"0057" => dat <= x"1283";
			when x"0058" => dat <= x"1303";
			when x"0059" => dat <= x"00A7";
			when x"005A" => dat <= x"1283";
			when x"005B" => dat <= x"1703";
			when x"005C" => dat <= x"0811";
			when x"005D" => dat <= x"3E15";
			when x"005E" => dat <= x"1783";
			when x"005F" => dat <= x"0084";
			when x"0060" => dat <= x"0800";
			when x"0061" => dat <= x"00D5";
			when x"0062" => dat <= x"1283";
			when x"0063" => dat <= x"1303";
			when x"0064" => dat <= x"1283";
			when x"0065" => dat <= x"1703";
			when x"0066" => dat <= x"0855";
			when x"0067" => dat <= x"1283";
			when x"0068" => dat <= x"1303";
			when x"0069" => dat <= x"00A7";
			when x"006A" => dat <= x"1283";
			when x"006B" => dat <= x"1703";
			when x"006C" => dat <= x"3001";
			when x"006D" => dat <= x"0791";
			when x"006E" => dat <= x"1803";
			when x"006F" => dat <= x"0A92";
			when x"0070" => dat <= x"3000";
			when x"0071" => dat <= x"0792";
			when x"0072" => dat <= x"0814";
			when x"0073" => dat <= x"3A80";
			when x"0074" => dat <= x"00D5";
			when x"0075" => dat <= x"0812";
			when x"0076" => dat <= x"3A80";
			when x"0077" => dat <= x"0255";
			when x"0078" => dat <= x"1D03";
			when x"0079" => dat <= x"287C";
			when x"007A" => dat <= x"0811";
			when x"007B" => dat <= x"0213";
			when x"007C" => dat <= x"1803";
			when x"007D" => dat <= x"287F";
			when x"007E" => dat <= x"2880";
			when x"007F" => dat <= x"2850";
			when x"0080" => dat <= x"0813";
			when x"0081" => dat <= x"00D5";
			when x"0082" => dat <= x"1283";
			when x"0083" => dat <= x"1303";
			when x"0084" => dat <= x"1283";
			when x"0085" => dat <= x"1703";
			when x"0086" => dat <= x"0855";
			when x"0087" => dat <= x"1283";
			when x"0088" => dat <= x"1303";
			when x"0089" => dat <= x"00A7";
			when x"008A" => dat <= x"1283";
			when x"008B" => dat <= x"1703";
			when x"008C" => dat <= x"0814";
			when x"008D" => dat <= x"01D7";
			when x"008E" => dat <= x"07D7";
			when x"008F" => dat <= x"0813";
			when x"0090" => dat <= x"01D6";
			when x"0091" => dat <= x"07D6";
			when x"0092" => dat <= x"3015";
			when x"0093" => dat <= x"120A";
			when x"0094" => dat <= x"118A";
			when x"0095" => dat <= x"2771";
			when x"0096" => dat <= x"120A";
			when x"0097" => dat <= x"118A";
			when x"0098" => dat <= x"2898";
			when x"0099" => dat <= x"2830";
			when x"009A" => dat <= x"120A";
			when x"009B" => dat <= x"118A";
			when x"009C" => dat <= x"2800";
			when x"0720" => dat <= x"00D8";
			when x"0721" => dat <= x"3000";
			when x"0722" => dat <= x"00D9";
			when x"0723" => dat <= x"3000";
			when x"0724" => dat <= x"00DA";
			when x"0725" => dat <= x"1003";
			when x"0726" => dat <= x"1283";
			when x"0727" => dat <= x"1303";
			when x"0728" => dat <= x"3000";
			when x"0729" => dat <= x"1803";
			when x"072A" => dat <= x"3001";
			when x"072B" => dat <= x"00A6";
			when x"072C" => dat <= x"0825";
			when x"072D" => dat <= x"1283";
			when x"072E" => dat <= x"1703";
			when x"072F" => dat <= x"00DB";
			when x"0730" => dat <= x"0859";
			when x"0731" => dat <= x"0758";
			when x"0732" => dat <= x"1783";
			when x"0733" => dat <= x"0084";
			when x"0734" => dat <= x"085B";
			when x"0735" => dat <= x"0080";
			when x"0736" => dat <= x"0859";
			when x"0737" => dat <= x"0758";
			when x"0738" => dat <= x"0084";
			when x"0739" => dat <= x"0800";
			when x"073A" => dat <= x"00DB";
			when x"073B" => dat <= x"1283";
			when x"073C" => dat <= x"1303";
			when x"073D" => dat <= x"1283";
			when x"073E" => dat <= x"1703";
			when x"073F" => dat <= x"085B";
			when x"0740" => dat <= x"1283";
			when x"0741" => dat <= x"1303";
			when x"0742" => dat <= x"00A7";
			when x"0743" => dat <= x"1283";
			when x"0744" => dat <= x"1703";
			when x"0745" => dat <= x"3001";
			when x"0746" => dat <= x"07D9";
			when x"0747" => dat <= x"1803";
			when x"0748" => dat <= x"0ADA";
			when x"0749" => dat <= x"3000";
			when x"074A" => dat <= x"07DA";
			when x"074B" => dat <= x"0859";
			when x"074C" => dat <= x"00DB";
			when x"074D" => dat <= x"1283";
			when x"074E" => dat <= x"1303";
			when x"074F" => dat <= x"1283";
			when x"0750" => dat <= x"1703";
			when x"0751" => dat <= x"085B";
			when x"0752" => dat <= x"1283";
			when x"0753" => dat <= x"1303";
			when x"0754" => dat <= x"00A7";
			when x"0755" => dat <= x"1283";
			when x"0756" => dat <= x"1703";
			when x"0757" => dat <= x"0859";
			when x"0758" => dat <= x"00DB";
			when x"0759" => dat <= x"1283";
			when x"075A" => dat <= x"1303";
			when x"075B" => dat <= x"1283";
			when x"075C" => dat <= x"1703";
			when x"075D" => dat <= x"085B";
			when x"075E" => dat <= x"1283";
			when x"075F" => dat <= x"1303";
			when x"0760" => dat <= x"00A6";
			when x"0761" => dat <= x"0825";
			when x"0762" => dat <= x"3A0A";
			when x"0763" => dat <= x"1D03";
			when x"0764" => dat <= x"2F66";
			when x"0765" => dat <= x"2F67";
			when x"0766" => dat <= x"2F2C";
			when x"0767" => dat <= x"1283";
			when x"0768" => dat <= x"1703";
			when x"0769" => dat <= x"085A";
			when x"076A" => dat <= x"01D7";
			when x"076B" => dat <= x"07D7";
			when x"076C" => dat <= x"0859";
			when x"076D" => dat <= x"01D6";
			when x"076E" => dat <= x"07D6";
			when x"076F" => dat <= x"2F70";
			when x"0770" => dat <= x"0008";
			when x"0771" => dat <= x"00D8";
			when x"0772" => dat <= x"3000";
			when x"0773" => dat <= x"00DA";
			when x"0774" => dat <= x"3000";
			when x"0775" => dat <= x"00DB";
			when x"0776" => dat <= x"3001";
			when x"0777" => dat <= x"00DC";
			when x"0778" => dat <= x"3000";
			when x"0779" => dat <= x"00DD";
			when x"077A" => dat <= x"2FDF";
			when x"077B" => dat <= x"1283";
			when x"077C" => dat <= x"1303";
			when x"077D" => dat <= x"0823";
			when x"077E" => dat <= x"3940";
			when x"077F" => dat <= x"1283";
			when x"0780" => dat <= x"1703";
			when x"0781" => dat <= x"00D9";
			when x"0782" => dat <= x"0859";
			when x"0783" => dat <= x"3A40";
			when x"0784" => dat <= x"1D03";
			when x"0785" => dat <= x"2F87";
			when x"0786" => dat <= x"2F88";
			when x"0787" => dat <= x"2FCC";
			when x"0788" => dat <= x"3001";
			when x"0789" => dat <= x"065C";
			when x"078A" => dat <= x"045D";
			when x"078B" => dat <= x"1D03";
			when x"078C" => dat <= x"2F8E";
			when x"078D" => dat <= x"2F8F";
			when x"078E" => dat <= x"2FAB";
			when x"078F" => dat <= x"3000";
			when x"0790" => dat <= x"00DC";
			when x"0791" => dat <= x"3000";
			when x"0792" => dat <= x"00DD";
			when x"0793" => dat <= x"085A";
			when x"0794" => dat <= x"0758";
			when x"0795" => dat <= x"1783";
			when x"0796" => dat <= x"0084";
			when x"0797" => dat <= x"0800";
			when x"0798" => dat <= x"00DE";
			when x"0799" => dat <= x"1283";
			when x"079A" => dat <= x"1303";
			when x"079B" => dat <= x"1283";
			when x"079C" => dat <= x"1703";
			when x"079D" => dat <= x"085E";
			when x"079E" => dat <= x"1283";
			when x"079F" => dat <= x"1303";
			when x"07A0" => dat <= x"00B8";
			when x"07A1" => dat <= x"16A4";
			when x"07A2" => dat <= x"1283";
			when x"07A3" => dat <= x"1703";
			when x"07A4" => dat <= x"3001";
			when x"07A5" => dat <= x"07DA";
			when x"07A6" => dat <= x"1803";
			when x"07A7" => dat <= x"0ADB";
			when x"07A8" => dat <= x"3000";
			when x"07A9" => dat <= x"07DB";
			when x"07AA" => dat <= x"2FCB";
			when x"07AB" => dat <= x"3002";
			when x"07AC" => dat <= x"065C";
			when x"07AD" => dat <= x"045D";
			when x"07AE" => dat <= x"1D03";
			when x"07AF" => dat <= x"2FB1";
			when x"07B0" => dat <= x"2FB2";
			when x"07B1" => dat <= x"2FCB";
			when x"07B2" => dat <= x"0857";
			when x"07B3" => dat <= x"065B";
			when x"07B4" => dat <= x"1D03";
			when x"07B5" => dat <= x"2FB8";
			when x"07B6" => dat <= x"0856";
			when x"07B7" => dat <= x"065A";
			when x"07B8" => dat <= x"1D03";
			when x"07B9" => dat <= x"2FBB";
			when x"07BA" => dat <= x"2FBC";
			when x"07BB" => dat <= x"2FC7";
			when x"07BC" => dat <= x"30DF";
			when x"07BD" => dat <= x"00DE";
			when x"07BE" => dat <= x"1283";
			when x"07BF" => dat <= x"1303";
			when x"07C0" => dat <= x"1283";
			when x"07C1" => dat <= x"1703";
			when x"07C2" => dat <= x"085E";
			when x"07C3" => dat <= x"1283";
			when x"07C4" => dat <= x"1303";
			when x"07C5" => dat <= x"05A4";
			when x"07C6" => dat <= x"2FCB";
			when x"07C7" => dat <= x"3001";
			when x"07C8" => dat <= x"00DC";
			when x"07C9" => dat <= x"3000";
			when x"07CA" => dat <= x"00DD";
			when x"07CB" => dat <= x"2FDF";
			when x"07CC" => dat <= x"08D9";
			when x"07CD" => dat <= x"1D03";
			when x"07CE" => dat <= x"2FD0";
			when x"07CF" => dat <= x"2FD1";
			when x"07D0" => dat <= x"2FDF";
			when x"07D1" => dat <= x"3002";
			when x"07D2" => dat <= x"00DC";
			when x"07D3" => dat <= x"3000";
			when x"07D4" => dat <= x"00DD";
			when x"07D5" => dat <= x"30DF";
			when x"07D6" => dat <= x"00DE";
			when x"07D7" => dat <= x"1283";
			when x"07D8" => dat <= x"1303";
			when x"07D9" => dat <= x"1283";
			when x"07DA" => dat <= x"1703";
			when x"07DB" => dat <= x"085E";
			when x"07DC" => dat <= x"1283";
			when x"07DD" => dat <= x"1303";
			when x"07DE" => dat <= x"05A4";
			when x"07DF" => dat <= x"1283";
			when x"07E0" => dat <= x"1703";
			when x"07E1" => dat <= x"0857";
			when x"07E2" => dat <= x"3A80";
			when x"07E3" => dat <= x"00DE";
			when x"07E4" => dat <= x"085B";
			when x"07E5" => dat <= x"3A80";
			when x"07E6" => dat <= x"025E";
			when x"07E7" => dat <= x"1D03";
			when x"07E8" => dat <= x"2FEB";
			when x"07E9" => dat <= x"085A";
			when x"07EA" => dat <= x"0256";
			when x"07EB" => dat <= x"1803";
			when x"07EC" => dat <= x"2FEE";
			when x"07ED" => dat <= x"2FEF";
			when x"07EE" => dat <= x"2F7B";
			when x"07EF" => dat <= x"085A";
			when x"07F0" => dat <= x"00DE";
			when x"07F1" => dat <= x"1283";
			when x"07F2" => dat <= x"1303";
			when x"07F3" => dat <= x"1283";
			when x"07F4" => dat <= x"1703";
			when x"07F5" => dat <= x"085E";
			when x"07F6" => dat <= x"1283";
			when x"07F7" => dat <= x"1303";
			when x"07F8" => dat <= x"00A7";
			when x"07F9" => dat <= x"3001";
			when x"07FA" => dat <= x"1283";
			when x"07FB" => dat <= x"1703";
			when x"07FC" => dat <= x"00DC";
			when x"07FD" => dat <= x"3000";
			when x"07FE" => dat <= x"00DD";
			when x"07FF" => dat <= x"0008";
			when x"2007" => dat <= x"3F72";
			when others => dat <= x"ffff";
		end case;
	end process;
end Behavioral;
